module adder (
	// inputs

	// outputs

);

endmodule


module top (
	// inputs

	// outputs

);


endmodule
